library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
entity control_memory is
port(
    MW : out std_logic;
    MM : out std_logic;
    RW : out std_logic;
    MD : out std_logic;
    FS : out std_logic_vector(4 downto 0);
    MB : out std_logic;
    TB : out std_logic;
    TA : out std_logic;
    TD : out std_logic;
    PL : out std_logic;
    PI : out std_logic;
    IL : out std_logic;
    MC : out std_logic;
    MS : out std_logic_vector(2 downto 0);
    NA : out std_logic_vector(7 downto 0);
    input : in std_logic_vector(7 downto 0);
    output : out std_logic_vector(27 downto 0)
);
end control_memory;
architecture behavioral of control_memory is
type mem_array is array(0 to 255) of std_logic_vector(27 downto 0);
begin
memory_m: process(input)
variable control_mem : mem_array:=(
    -- 0
    x"C020224", -- 0    ADI
    x"C02000C", -- 1    LD
    x"C020001", -- 2    ST 
    x"C020014", -- 3    INC
    x"C0200E4", -- 4    NOT
    x"C020024", -- 5    ADD
    x"C022000", -- 6    B
    x"C880000", -- 7    BZ
    x"C020000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- 1
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- 2
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- 3
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- 4
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- 5
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- 6
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- 7
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- 8
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- 9
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- A
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- B
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- C
    x"C100002", -- 0
    x"C20C002", -- 1
    x"0030000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"C022000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- D
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- E
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000", -- F
    -- F
    x"0000000", -- 0
    x"0000000", -- 1
    x"0000000", -- 2
    x"0000000", -- 3
    x"0000000", -- 4
    x"0000000", -- 5
    x"0000000", -- 6
    x"0000000", -- 7
    x"0000000", -- 8
    x"0000000", -- 9
    x"0000000", -- A
    x"0000000", -- B
    x"0000000", -- C
    x"0000000", -- D
    x"0000000", -- E
    x"0000000" -- F
);
variable address : integer;
variable control_out : std_logic_vector(27 downto 0);
begin
    address := conv_integer(input);
    control_out := control_mem(address);
    output <= control_out;
    MW <= control_out(0);
    MM <= control_out(1);
    RW <= control_out(2);
    MD <= control_out(3);
    FS <= control_out(8 downto 4);
    MB <= control_out(9);
    TB <= control_out(10);
    TA <= control_out(11);
    TD <= control_out(12);
    PL <= control_out(13);
    PI <= control_out(14);
    IL <= control_out(15);
    MC <= control_out(16);
    MS <= control_out(19 downto 17);
    NA <= control_out(27 downto 20);
end process;
end behavioral;
